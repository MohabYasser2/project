
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY MEMORY IS

PORT (
CLK,RST,PUSH,POP,MEM_WRITE,INTERRUPT_SIG,MEMTOREG:IN std_logic;
ALU_OUTPUT: IN std_logic_vector(31 DOWNTO 0);
Write_DATA: IN std_logic_vector(31 DOWNTO 0);
MEM_OUTPUT: OUT  std_logic_vector(31 DOWNTO 0);
FLAGS: IN std_logic_vector(3 downto 0);
BRANCH_SIG_IN : IN std_logic;
BRANCH_Z_SIG_IN : IN std_logic;
Protect_sig : IN std_logic;
Free_sig: IN STD_LOGIC;
PC: IN std_logic_vector(31 DOWNTO 0);
callSig: IN STD_LOGIC;
RET_SIG: IN STD_LOGIC;
RTI_SIG: IN STD_LOGIC;

RET_SIG_OUT: OUT STD_LOGIC;
RTI_SIG_OUT: OUT STD_LOGIC;
BRANCH_SIG : OUT std_logic;
BRANCH_Z_SIG : OUT std_logic;
FLUSH_SIG: OUT STD_LOGIC;
Flags_out: OUT std_logic_vector(3 DOWNTO 0);

EXCEPTION_O : OUT STD_LOGIC
);

END ENTITY;

Architecture FetchUnit of MEMORY IS

component INC_DEC IS
PORT(	CLK, RST,PUSH,POP,CALL_SIG,RET_SIG,RTI_SIG,INTERRUPT_SIG: IN STD_LOGIC;
DATAIN: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
DATAOUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END component;

component SP IS
	PORT(	CLK, RST: IN STD_LOGIC;
		DATAIN: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATAOUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END component;

Component DataMemory IS

PORT (
CLK,RST,WE,INTERRUPT_SIG,RTI_SIG,MEMTOREG: IN std_logic;
Protect_SIG,Free_SIG : IN std_logic;
ADDRESS : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
WriteData: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
FLAGS: IN STD_LOGIC_VECTOR(3 DOWNTO 0):= (OTHERS => '0');
DATAOUT : OUT std_logic_vector(31 DOWNTO 0);
FLAGS_OUT: OUT std_logic_vector(3 DOWNTO 0);
EXCEPTION_OUT : OUT STD_LOGIC
);

END component;

component Mux2x1 IS
generic(N : INTEGER );
PORT(
I0,I1: IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
S : IN STD_LOGIC;
O : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0 ));

END component;

--Signals
Signal MUXOUT : std_logic_vector(31 DOWNTO 0);
Signal SP_TEMP : std_logic_vector(31 downto 0);
Signal INC_DEC_OUTPUT : std_logic_vector(31 downto 0);
signal OR_OUTPUT,OR_OUTPUT2 : std_logic;
Signal Dout : std_logic_vector(31 DOWNTO 0);
--Signal FLAGS_OUT : std_logic_vector(3 DOWNTO 0); --USE IN RTI


BEGIN
OR_OUTPUT <= POP OR PUSH OR CallSIG OR RET_SIG OR RTI_SIG OR INTERRUPT_SIG;
OR_OUTPUT2 <= CallSIG OR INTERRUPT_SIG;
BRANCH_SIG <= BRANCH_SIG_IN;

BRANCH_Z_SIG <= BRANCH_Z_SIG_IN AND FLAGS(0);

FLUSH_SIG <= CALLSIG OR RET_SIG OR RTI_SIG OR INTERRUPT_SIG;
RET_SIG_OUT <= RET_SIG;
RTI_SIG_OUT <= RTI_SIG;


U0:Mux2x1 GENERIC MAP (32) PORT MAP(ALU_OUTPUT,SP_TEMP ,OR_OUTPUT,MUXOUT);

U4:Mux2x1 GENERIC MAP (32) PORT MAP(Write_data,PC ,OR_OUTPUT2,Dout);

U1:DATAMEMORY PORT MAP(CLK,RST,MEM_WRITE,INTERRUPT_SIG,RTI_SIG,MEMTOREG,Protect_SIG,Free_Sig,MUXOUT,Dout,FLAGS,MEM_OUTPUT,FLAGS_OUT,EXCEPTION_O);

U2:SP Port MAP(CLK,RST,INC_DEC_OUTPUT,SP_TEMP);

U3:INC_DEC Port MAP(CLK,RST,PUSH,POP,Callsig,RET_SIG,RTI_SIG,INTERRUPT_SIG,SP_TEMP,INC_DEC_OUTPUT);


END ARCHITECTURE;