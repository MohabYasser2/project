LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CCR IS
	PORT(
		CLK, RST,RTI_SIG : IN STD_LOGIC;
		DATAIN: IN STD_LOGIC_VECTOR(3 downto 0);
		RTI_FLAGS: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATAOUT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE CCR_ARCH OF CCR IS
	SIGNAL DATA: STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
BEGIN
	PROCESS(CLK, RST) IS
	
	BEGIN
		IF RST = '1' THEN
			DATA<= (OTHERS => '0');
		ELSIF RISING_EDGE(CLK)  THEN
			IF RTI_SIG = '1' THEN
				DATA <= RTI_FLAGS;
			ELSE
				DATA <= STD_LOGIC_VECTOR(UNSIGNED(DATAIN));
			END IF;
		END IF;
	END PROCESS;
	DATAOUT<= DATA ;
	
	END ARCHITECTURE;
