LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY REGISTERFILE32 IS

PORT (
CLK, RST, WE : IN std_logic;
DATAIN : IN std_logic_vector(31 DOWNTO 0);
READADDRESS1, READADDRESS2, WRITEADDRESS : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
DATAOUT1, DATAOUT2 : OUT std_logic_vector(31 DOWNTO 0)
);

END ENTITY;

ARCHITECTURE ARCH OF REGISTERFILE32 IS

TYPE ram_type IS ARRAY(7 DOWNTO 0) of std_logic_vector(31 DOWNTO 0);
SIGNAL RAM : ram_type ;

BEGIN

PROCESS(CLK, RST) IS
BEGIN

IF RST = '1' THEN

RAM <= (OTHERS => (OTHERS => '0'));

ELSIF falling_edge(CLK) THEN
IF WE = '1' THEN
RAM(to_integer(unsigned(WRITEADDRESS))) <= DATAIN;
END IF;
END IF;

END PROCESS;

DATAOUT1 <= RAM(to_integer(unsigned(READADDRESS1)));
DATAOUT2 <= RAM(to_integer(unsigned(READADDRESS2)));

END ARCHITECTURE;
