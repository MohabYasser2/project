
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY M_WB IS
	PORT(	CLK, RST: IN STD_LOGIC;
		MemToReg,RegWrite,In_SIG: IN STD_LOGIC;
		MEM_OUTPUT,ALU_OUTPUT,IN_PORT: IN STD_LOGIC_VECTOR(31 DOWNTO 0); 
		Write_Address: IN STD_LOGIC_VECTOR(2 DOWNTO 0); 
		SWAPPING: IN STD_LOGIC;
		MemToReg_OUT,RegWrite_OUT,In_SIG_OUT: OUT STD_LOGIC;
		MEM_OUTPUT_OUT,ALU_OUTPUT_OUT,IN_PORT_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0); 
		Write_Address_OUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		SWAPPING_OUT: OUT STD_LOGIC





);
		
END ENTITY;

ARCHITECTURE FDREGARCH OF M_WB IS
BEGIN

	PROCESS(CLK) IS
	BEGIN
		
		IF RISING_EDGE(CLK) THEN

			IF RST = '1' THEN
			MemToReg_OUT <= '0';
			RegWrite_OUT <= '0';
			In_SIG_OUT <= '0';
			MEM_OUTPUT_OUT  <= (OTHERS => '0');
			ALU_OUTPUT_OUT <= (OTHERS => '0');
			IN_PORT_OUT <= (OTHERS => '0');
			Write_Address_OUT <= (OTHERS => '0');
			SWAPPING_OUT <= '0';
			ELSE
			MemToReg_OUT <= MemToReg;
			RegWrite_OUT <= RegWrite;
			In_SIG_OUT <= In_SIG;
			MEM_OUTPUT_OUT  <= MEM_OUTPUT;
			ALU_OUTPUT_OUT <= ALU_OUTPUT;
			IN_PORT_OUT <= IN_PORT;
			Write_Address_OUT <= Write_Address;
			SWAPPING_OUT <= SWAPPING;
			END IF; 

		END IF;
	END PROCESS;

END ARCHITECTURE;



