LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY INSTRUCTION_CACHE IS

PORT (
CLK, RST : IN std_logic;
PC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
DATAOUT : OUT std_logic_vector(15 DOWNTO 0);
RESET_VALUE : OUT std_logic_vector(31 DOWNTO 0)

);

END ENTITY;

ARCHITECTURE ARCH OF INSTRUCTION_CACHE IS
signal DATA : std_logic_vector(15 DOWNTO 0);
TYPE ram_type IS ARRAY(4095 DOWNTO 0) of std_logic_vector(15 DOWNTO 0);
SIGNAL INSTRUCTION_CACHE : ram_type ;

BEGIN

PROCESS(RST,CLK) IS
BEGIN

IF RST = '1' THEN

INSTRUCTION_CACHE <= (OTHERS => (OTHERS => '0'));

END IF;

IF FALLING_EDGE(CLK) THEN
DATA <=INSTRUCTION_CACHE(to_integer(unsigned(PC)));
END IF;

END PROCESS;

DATAOUT <= DATA;
RESET_VALUE <= INSTRUCTION_CACHE(1) & INSTRUCTION_CACHE(0);

END ARCHITECTURE;
