
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SP IS
	PORT(	CLK, RST: IN STD_LOGIC;
		DATAIN: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATAOUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE SP_ARCH OF SP IS
	

	SIGNAL TEMP_DATAIN: STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000011111111111" ;
BEGIN
	PROCESS(CLK, RST) IS
	
	BEGIN
		IF RST = '1' THEN
			Temp_DATAIN <= "00000000000000000000011111111111";
		ELSIF RISING_EDGE(CLK) 
		THEN
			Temp_DATAIN <= DATAIN;
		END IF;
	END PROCESS;
	
	DATAOUT <= Temp_DATAIN;

END ARCHITECTURE;